"Mon Mar 12 15:06:50 CET 2018";"@Teranga News";"New";"post:";"Phase";"II";"du";"PUDC";":";"Souleymane";"Jules";"Diop";"annonce";"la";"https://t.co/KenMFyBk5K";"#Fatick";"#NEPAD";"#PUDC";"#CESTMOB";"#kebetu";"#Senegal"
"Mon Mar 12 15:06:23 CET 2018";"@Sophie Ndiaye Sy";"RT";"@imajeader:";"Le";"Super";"Women";"Leadership";"Conference";"2018";"de";"JEADER";"SENEGAL,";"ce";"sera";"ce";"Samedi";"17";"au";"Novotel";"sous";"le";"thème";"de";"la";"Trans'Missi…"
"Mon Mar 12 15:06:04 CET 2018";"@Hayssatu";"RT";"@SySeynabou:";"J'invite";"mes";"amis,chercheurs";"ou";"pas,";"qui";"se";"sentent";"concernés";"de";"constituer";"une";"équipe";"pluridisciplinaire";"et";"faire";"1";"étude…"
"Mon Mar 12 15:05:43 CET 2018";"@finance news Turkey";"RT";"@MevlutCavusoglu:";"#Türkiye-#Senegal";"işbirliği";"meyvelerini";"veriyor,";"ekonomik";"ve";"ticari";"ilişkilerde";"hedefler";"aşılıyor.";"İkili";"ticaret";"hacmi…"
"Mon Mar 12 15:05:38 CET 2018";"@Jummy Thompson";"RT";"@NaijaBet:";"Today's";"Fixtures";"⚽";"";"England-";"Premier";"League";"2";"International";"Youth-";"Viareggio";"Youth";"Cup";"Senegal-";"Premier";"League";"Belgium-";"U21,…"
"Mon Mar 12 15:05:27 CET 2018";"@Didier vevo";"RT";"@Cherif221:";""Un";"véhicule";"de";"gendarmes";"(avec";"des";"détenus)";"qui";"roule";"en";"sens";"inverse";"sur";"une";"bretelle";"de";"l’autoroute.";"Bien";"évidemment";"l’ir…"
"Mon Mar 12 15:05:23 CET 2018";"@SENY";"RT";"@apapanne:";"Wallah";"l'eau";"que";"nous";"donne";"la";"@senegal_SDE";"c'est";"une";"grosse";"farce.";"On";"dirait";"que";"tu";"prends";"un";"médicament.";"Respectez";"nous";"qua…"
"Mon Mar 12 15:05:12 CET 2018";"@United boy";"RT";"@statsgh:";"It";"is";"cheaper";"to";"travel";"by";"air";"from";"Accra";"to";"London";"than";"from";"Accra";"to";"Dakar";"(Senegal)";"which";"is";"in";"West";"Africa."
"Mon Mar 12 15:04:58 CET 2018";"@No one";"RT";"@SySeynabou:";"J'invite";"mes";"amis,chercheurs";"ou";"pas,";"qui";"se";"sentent";"concernés";"de";"constituer";"une";"équipe";"pluridisciplinaire";"et";"faire";"1";"étude…"
"Mon Mar 12 15:04:42 CET 2018";"@DakarFlash";"#Senegal";"Cheikh";"Traoré";":";"«";"Si";"Fada";"rejoint";"Macky,";"je";"le";"quitte";"sans";"réfléchir";"»";"https://t.co/cx7mwqLYKq"
"Mon Mar 12 15:04:23 CET 2018";"@senegal7";"Vidéo:";"Mamadou";"Faye,";"premier";"président";"de";"la";"cour";"des";"comptes:";""Ce";"que";"nous";"déplorons,";"c'est..."";"-";"https://t.co/yG2Cyhcj60";"#Senegal";"#Kebetu";"#Dakar";"#team221";"#Mali";"#Mauritanie";"https://t.co/yuY6eJyL7F"
"Mon Mar 12 15:03:53 CET 2018";"@ILOVESENEGAL";"RT";"@Marie88838201:";"@KeryJames";"Le";"Sénégal";"🇸🇳";"🙏🏼♥️"
"Mon Mar 12 15:03:08 CET 2018";"@koaci.com";"Sénégal:";"Akon";"candidat";"Présidentielle";"américaine";"de";"2020";"Mark";"Zuckerberg";"comme";"colistier...";"https://t.co/0Ny68IesKT"
"Mon Mar 12 15:03:02 CET 2018";"@Fall Mambaye";"RT";"@hadyba_:";"On";"dirait";"que";"le";"Sénégal";"a";"son";"BHL.";"Je";"connais";"M.";"Diouf.";"On";"collaborait";"jusqu'à";"cette";"année";"dans";"l'encadrement";"des";"stagiaires.…"
"Mon Mar 12 15:02:55 CET 2018";"@SeneNews";"Népal:";"";"prés";"de";"40";"morts";"enregistrés";"dans";"un";"crash";"d’avion";"à";"l’aéroport";"de";"Katmandou";"#kebetu";"#senegal";"https://t.co/2XQ26iUBxf";"https://t.co/rlPXcKubAv"
"Mon Mar 12 15:02:48 CET 2018";"@wiwsport.com";"Keita";"Baldé";"et";"Ferland";"Mendy";"dans";"l'équipe";"type";"de";"la";"29e";"journée";"de";"Ligue";"1";"#Senegal";"#wiwsport";">";"https://t.co/oH84RQA1Ly";"https://t.co/LD7JLy7xuv";"https://t.co/hrL4NNSaGS"
"Mon Mar 12 15:02:30 CET 2018";"@koaci.com";"Sénégal:";"Akon";"candidat";"Présidentielle";"américaine";"de";"2020";"Mark";"Zuckerberg";"comme";"colistier";"https://t.co/wyvuFnimmi"
"Mon Mar 12 15:02:28 CET 2018";"@Barrow-Meter";"RT";"@BarrowPresident:";"We";"belief";"in";"strengthening";"bilateral";"ties";"for";"the";"socio-economic";"and";"political";"benefits";"of";"our";"people.";"";"I";"am";"honoured…"
"Mon Mar 12 15:02:20 CET 2018";"@J. Lawal #IBLFellow";"RT";"@ABANAngels:";"Senegal's";"recent";"30-year";"$1";"billion";"Eurobond";"attracted";"a";"coupon";"rate";"of";"6.75%";"-";"the";"lowest";"among";"other";"recent";"African";"issue…"
"Mon Mar 12 15:02:18 CET 2018";"@Inspecteurgadget";"RT";"@__Diarra:";"Gniy";"participer";"si";"#";"bi";"pour";"Sénégal,";"douggeul";"lène";"vos";"beaux";"yéré";"wolof";"way";"ngey";"représenter";"culture";"bi"
"Mon Mar 12 15:02:14 CET 2018";"@Rene Lake";"Tant";"pis";"si";"certains";"Sénégalais";"n’aiment";"pas";"les";"bonnes";"nouvelles,";"mais";"de";"bonnes";"performances";"économiques,";"la";"gouvernance";"du";"Président";"#Macky";"Sall";"en";"a";"réalisé";"";"-";"L’opposition";"préfère";"détourner";"le";"regard";"et";"se";"boucher";"les";"oreilles.";"#Kebetu";"#Sénégal";"➡https://t.co/MC4XQA0vSC";"https://t.co/qtJ3EVoOUB"
"Mon Mar 12 15:02:14 CET 2018";"@SenePlus.com";"Tant";"pis";"si";"certains";"Sénégalais";"n’aiment";"pas";"les";"bonnes";"nouvelles,";"mais";"de";"bonnes";"performances";"économiques,";"la";"gouvernance";"du";"Président";"#Macky";"Sall";"en";"a";"réalisé";"";"-";"L’opposition";"préfère";"détourner";"le";"regard";"et";"se";"boucher";"les";"oreilles.";"#Kebetu";"#Sénégal";"➡https://t.co/MPeg75ZsH1";"https://t.co/7HuWlJjRuq"
"Mon Mar 12 15:01:42 CET 2018";"@Ubuntu Africa Chile";"@PapinoMatus";"siguenos,";"pronto";"tenemos";"la";"fiesta";"de";"senegal";"el";"7";"de";"abril"
"Mon Mar 12 15:01:35 CET 2018";"@Ney Ney 🇸🇳⚡️";"RT";"@BaalbakiFootbal:";"@SenegalFootball";"@Macky_Sall";"@PR_Senegal";"Nos";"lions";"nous";"ont";"fait";"rêver";"en";"2002";"pour";"atteindre";"les";"1/4";"F";"de";"la";"coupe";"du…"
"Mon Mar 12 15:01:23 CET 2018";"@Shaykh Ibraheem";"Wallah";"l'eau";"que";"nous";"donne";"la";"@senegal_SDE";"c'est";"une";"grosse";"farce.";"On";"dirait";"que";"tu";"prends";"un";"médicament.";"Respectez";"nous";"quand";"même"
"Mon Mar 12 15:01:21 CET 2018";"@Rachel Léa";"RT";"@SySeynabou:";"J'invite";"mes";"amis,chercheurs";"ou";"pas,";"qui";"se";"sentent";"concernés";"de";"constituer";"une";"équipe";"pluridisciplinaire";"et";"faire";"1";"étude…"
"Mon Mar 12 15:00:44 CET 2018";"@Queen Things Podcast";"#Senegal";"#America";"-";"@issarae";"is";"an";"actress,";"writer,";"director,";"producer,";"and web";"series creator.";"She";"first";"attracted";"attention";"for";"her";"work";"on";"the YouTube web";"series Awkward";"Black";"Girl";"and HBO television";"series Insecure";"#QueenThingsOnly";"#AfricanQueensProject";"https://t.co/JZR3TGYxlt"
"Mon Mar 12 15:00:36 CET 2018";"@Nopiwouma";"RT";"@SySeynabou:";"J'invite";"mes";"amis,chercheurs";"ou";"pas,";"qui";"se";"sentent";"concernés";"de";"constituer";"une";"équipe";"pluridisciplinaire";"et";"faire";"1";"étude…"
"Mon Mar 12 15:00:33 CET 2018";"@Dagnogo Naga Inza";"RT";"@SySeynabou:";"J'invite";"mes";"amis,chercheurs";"ou";"pas,";"qui";"se";"sentent";"concernés";"de";"constituer";"une";"équipe";"pluridisciplinaire";"et";"faire";"1";"étude…"
"Mon Mar 12 15:00:25 CET 2018";"@Ondoua Akoa georges";"Avis";"d’appel";"d’offres";"ouvert";"à";"l’international";"au";"Sénégal";"https://t.co/GSuVCajuu1";"https://t.co/aO9KVqhdVj"
"Mon Mar 12 15:00:13 CET 2018";"@мoиzεя | مُنذّر ♕";"RT";"@_Mazin777:";"That’s";"it,";"I’m";"moving";"to";"senegal";"https://t.co/0ev4810pX5"
"Mon Mar 12 15:00:10 CET 2018";"@DakarFlash";"#Senegal";"Discours";"de";"Sidy";"Lamine";"Niasse";":";"une";"attaque";"en";"règle";"contre";"son";"frère";"l’imam";"Araby";"Niasse";"?";"https://t.co/Bwq3yxiN7n"
"Mon Mar 12 15:00:05 CET 2018";"@senegalbot";"RT";"@teledakar:";"#kebetu";"#senegal";"Vous";"cherchez";"des";"visas";":";"Évitez";"ces";"deux";"femmes...";"Regardez";"!";"https://t.co/AlBgVBpd6K"
"Mon Mar 12 15:00:05 CET 2018";"@senegalbot";"RT";"@cuisineanxious:";"Alors";"qu'il";"n'a";"que";"10";"ans,";"le";"père";"de";"Camille";"Millerand";"l’emmène";"en";"Afrique";"(un";"continent";"qu'il";"ne";"connait";"pas).";"Ils";"p…"
"Mon Mar 12 15:00:05 CET 2018";"@senegalbot";"RT";"@RIBETTAR:";"Idrissa";"Seck";":";"«";"La";"première";"maladie";"du";"Sénégal,";"c’est";"Macky";"Sall";"»";"https://t.co/RtkNRWNkb3";"on";"@bloglovin"
"Mon Mar 12 15:00:05 CET 2018";"@aDakar";"#Senegal";"Procédures";"de";"passation";"des";"marchés";"Le";"Coud";"démonte";"le";"rapport";"de";"l’ARMP";"#aDakar";"https://t.co/7HFqIkRc5C"
"Mon Mar 12 15:00:04 CET 2018";"@senegalbot";"RT";"@RIBETTAR:";"Le";"Sénégal";"extrade";"en";"Mauritanie";"un";"Français,";"trafiquant";"de";"drogue";"https://t.co/RgRK8ET1lj";"on";"@bloglovin"
"Mon Mar 12 15:00:04 CET 2018";"@senegalbot";"RT";"@XoromD:";"@AprChine";"@Macky_Sall";"@elhadjkasse";"@tallamouna";"@MosesSarr";"@PR_Senegal";"@aidadpeters";"@FayeSallMarieme";"@HashtagSenegaal";"@avecmacky…"
"Mon Mar 12 15:00:03 CET 2018";"@senegalbot";"RT";"@stopscammerscom:";"Romance";"Scammer:";"Basirat";"Ibrahim";"25";"y.o.";"from";"Dakar";"(Senegal)";"https://t.co/lzzBNvioTC"
"Mon Mar 12 15:00:03 CET 2018";"@FranceMondeNews";"Sénégal";":";"le";"combat";"des";"grandes";"sœurs";"contre";"l'excision";"https://t.co/l7bwiC7TaH";":Auto";"pickup";"by";"wikyou"
"Mon Mar 12 15:00:03 CET 2018";"@senegalbot";"RT";"@Nabou_shou:";"@khouma_racky";"";"take!";"So";"i’am";"too";"late";"#FinePeoplefromSenegal";"";"Senegal";"rek";"🌺💎";"https://t.co/HUHgaLvjdK"
"Mon Mar 12 15:00:03 CET 2018";"@senegalbot";"RT";"@Marsattaqueblog:";"Sur";"les";"+1.850";"postes";"dédiés";"aux";"unités";"opérationnelles";"et";"leur";"environnement";"sur";"la";"#LPM";"2019-2025";"(sur";"les";"6.000";"au…"
"Mon Mar 12 15:00:02 CET 2018";"@senegalbot";"RT";"@Pressafrik:";"Victoire";"de";"Boy";"Niang";"2";":";"«";"Moustapha";"Gueye";"a";"donné";"la";"clé";"qui";"battu";"Sa";"Thiès";"»,";"selon";"le";"père";"de";"Boye";"Niang";"2";"Ce";"dimanche,…"
"Mon Mar 12 15:00:02 CET 2018";"@senegalbot";"RT";"@IbrahimNdiaye9:";""Le";"système";"politique";"#Senegal-ais";"est";"électoralo-centriste",";"selon";"le";"professeur";"Jean-Charles";"Biagui.";"C'est";"dire";"que";"l…"
"Mon Mar 12 15:00:00 CET 2018";"@Befoune.";"RT";"@SySeynabou:";"J'invite";"mes";"amis,chercheurs";"ou";"pas,";"qui";"se";"sentent";"concernés";"de";"constituer";"une";"équipe";"pluridisciplinaire";"et";"faire";"1";"étude…"
"Mon Mar 12 14:59:47 CET 2018";"@Ibrahim Ndiaye";""Le";"système";"politique";"#Senegal-ais";"est";"électoralo-centriste",";"selon";"le";"professeur";"Jean-Charles";"Biagui.";"C'est";"dire";"que";"la";"démocratie";"ne";"résume";"pas";"qu'aux";"élections.";"#Senegal";"#Politique"
"Mon Mar 12 14:59:36 CET 2018";"@Cheick Oumar Diallo";"RT";"@yeesalagrihub:";"Que";"veut";"dire";"Yeesal";"?";"Yeesal";"est";"un";"terme";"wolof";"qui";"signifie";"“innover”";"ou";"“rénover”.";"Ce";"nom";"a";"été";"choisi";"pour";"se";"confor…"
"Mon Mar 12 14:59:21 CET 2018";"@DoroFineGirl";"RT";"@SySeynabou:";"J'invite";"mes";"amis,chercheurs";"ou";"pas,";"qui";"se";"sentent";"concernés";"de";"constituer";"une";"équipe";"pluridisciplinaire";"et";"faire";"1";"étude…"
"Mon Mar 12 14:59:16 CET 2018";"@CouscousBoulette";"RT";"@PR_Senegal:";"Le";"Chef";"de";"l’Etat";"@Macky_Sall";"a";"présidé";"hier";"la";"cérémonie";"officielle";"de";"présentation";"du";"#TrophyTour";"de";"la";"Coupe";"du";"monde";"de…"
"Mon Mar 12 14:58:56 CET 2018";"@Pressafrik.com";"Victoire";"de";"Boy";"Niang";"2";":";"«";"Moustapha";"Gueye";"a";"donné";"la";"clé";"qui";"battu";"Sa";"Thiès";"»,";"selon";"le";"père";"de";"Boye";"Niang";"2";"Ce";"dimanche,";"le";"combat";"Sa";"Thiès-Boy";"Niang";"2";"a";"tenu";"les";"férus";"de";"lutte.&nbsp;";"Le";"second";"nommé";"a";"battu";"en";"moins";"de";"deux...";"|";"#kebetu";"#Senegal";"https://t.co/HTfbHkGgXB";"https://t.co/YqKsKsSrCR"
"Mon Mar 12 14:58:53 CET 2018";"@Clé De La Réussite";"RT";"@KeryJames:";"Photo";"prise";"sur";"l'île";"de";"Gorée";"au";"#Senegal.";"https://t.co/TdOw6SJawK"
"Mon Mar 12 14:58:51 CET 2018";"@Santana M";"RT";"@nialaruh_:";"Yasss";"I’m";"moving";"to";"Senegal";"https://t.co/V4sDraG3Xj"
"Mon Mar 12 14:58:47 CET 2018";"@FdeStV";"Sur";"les";"+1.850";"postes";"dédiés";"aux";"unités";"opérationnelles";"et";"leur";"environnement";"sur";"la";"#LPM";"2019-2025";"(sur";"les";"6.000";"au";"total),";"environ";"300";"bénéficieront";"aux";"forces";"de";"présence";"et";"de";"souveraineté";"(notamment";"dans";"le";"soutien)";":";"Sénégal,";"Djibouti,";"Guyane,";"La";"Réunion,";"etc.";"#armées"
"Mon Mar 12 14:58:23 CET 2018";"@Mery";"RT";"@nopiwouma:";"On";"ne";"peut";"pas";"tolérer";"le";"genre";"de";"propos";"que";"le";"Pr";"Songué";"Diouf";"sur";"@tfm_senegal";"faisant";"l'apologie";"du";"viol!";"Protégez";"nos";"f…"
"Mon Mar 12 14:57:46 CET 2018";"@afrofeminista";"RT";"@SySeynabou:";"J'invite";"mes";"amis,chercheurs";"ou";"pas,";"qui";"se";"sentent";"concernés";"de";"constituer";"une";"équipe";"pluridisciplinaire";"et";"faire";"1";"étude…"
"Mon Mar 12 14:57:19 CET 2018";"@Nabou’shou🌺💎";"@khouma_racky";"";"take!";"So";"i’am";"too";"late";"#FinePeoplefromSenegal";"";"Senegal";"rek";"🌺💎";"https://t.co/HUHgaLvjdK"
"Mon Mar 12 14:57:03 CET 2018";"@Stop-Scammers.com";"Romance";"Scammer:";"Basirat";"Ibrahim";"25";"y.o.";"from";"Dakar";"(Senegal)";"https://t.co/lzzBNvioTC"
"Mon Mar 12 14:56:55 CET 2018";"@@.🇸🇳";"@AprChine";"@Macky_Sall";"@elhadjkasse";"@tallamouna";"@MosesSarr";"@PR_Senegal";"@aidadpeters";"@FayeSallMarieme";"@HashtagSenegaal";"@avecmackysall";"@AvecMacky";"@BBYSenegal";"@partageleen";"@LioMdX";"@amadoud98130314";"@djibrilsene24";"@darkologi";"@moussadiallovl";"@ThereseaidaS";"@cherif_aidara1";"@aissatousaneh";"@shaia_fall";"@KaneRaki";"@ado_cisse";"Je";"fais";"allusion";"à";"la";"France...";"puisse";"que";"c’";"est";"votre";"référence";".pas";"la";"présence";"de";"Macron";"ou";"d’";"un";"ministre.."
"Mon Mar 12 14:56:29 CET 2018";"@Collateral Beauty";"RT";"@Ares210:";"Je";"suis";"indigné";"et";"choqué";"par";"les";"propos";"diffusés";"par";"@tfm_senegal";"@GFMofficiel";"durant";"l'émission";"#JakaarloBi";"Ce";"discours";"est…"
"Mon Mar 12 14:56:29 CET 2018";"@Essongori Maribau";"RT";"@AmbaPikin:";"@_AfricanUnion";"should";"do";"the";"right";"thing";"and";"show";"the";"world";"it's";"not";"made";"up";"of";"#shitholecountries";"#SuspendCameroun";"Free";"#Am…"
"Mon Mar 12 14:56:27 CET 2018";"@Otunba (Engr.) MOOB";"RT";"@smallstarters:";"Meet";"the";"33-year-old";"lady";"at";"the";"helm";"of";"#Senegal's";"biggest";"poultry";"company";"";"https://t.co/N2qeM5slwk";"";"Anta";"Babacar";"Ngom…"
"Mon Mar 12 14:56:11 CET 2018";"@🎢";"RT";"@_therealbene:";"Continue";"à";"ne";"pas";"voir";"alors.";"Deja";"le";"prix";"du";"billet";"n'est";"pas";"le";"même";"que";"celui";"du";"Sénégal";"ou";"Mali,";"ensuite";"en";"ce";"moment…"
"Mon Mar 12 14:56:10 CET 2018";"@#MGWV ★ RIBETTAR";"Le";"Sénégal";"extrade";"en";"Mauritanie";"un";"Français,";"trafiquant";"de";"drogue";"https://t.co/RgRK8ET1lj";"on";"@bloglovin"
"Mon Mar 12 14:56:10 CET 2018";"@#MGWV ★ RIBETTAR";"Idrissa";"Seck";":";"«";"La";"première";"maladie";"du";"Sénégal,";"c’est";"Macky";"Sall";"»";"https://t.co/RtkNRWNkb3";"on";"@bloglovin"
"Mon Mar 12 14:56:08 CET 2018";"@Simon Decreuze";"Alors";"qu'il";"n'a";"que";"10";"ans,";"le";"père";"de";"Camille";"Millerand";"l’emmène";"en";"Afrique";"(un";"continent";"qu'il";"ne";"connait";"pas).";"Ils";"partent";"en";"camion";"et";"logent";"chez";"l'habitant";"et";"vont";"traverser";"le";"Maroc,";"la";"Mauritanie,";"le";"Sénégal,";"la";"Guinée";"Conakry";"et";"la";"Côte";"d'Ivoire...La";"suite";"est";"à";"écouter";"https://t.co/82BQ18UqzR"
"Mon Mar 12 14:56:06 CET 2018";"@Teledakar";"#kebetu";"#senegal";"Vous";"cherchez";"des";"visas";":";"Évitez";"ces";"deux";"femmes...";"Regardez";"!";"https://t.co/AlBgVBpd6K"
"Mon Mar 12 14:55:50 CET 2018";"@Claudia";"RT";"@RiscattoNaz:";"E";"per";"la";"madre";"di";"Pamela";"Mastropietro??";"https://t.co/V5kDcmvkaL";"via";"@RiscattoNaz"
"Mon Mar 12 14:55:43 CET 2018";"@Anne-Laure GRIMAUD";"RT";"@Ju_Alemany:";"L'aventure";"commence";"ici";"https://t.co/Ee1iDhoYy3";"https://t.co/Oj42wuR5aV"
"Mon Mar 12 14:55:14 CET 2018";"@Inspecteurgadget";"RT";"@PR_Senegal:";"Le";"Chef";"de";"l’Etat";"@Macky_Sall";"a";"présidé";"hier";"la";"cérémonie";"officielle";"de";"présentation";"du";"#TrophyTour";"de";"la";"Coupe";"du";"monde";"de…"
"Mon Mar 12 14:54:46 CET 2018";"@NFatou Kane ♐️🎀📚";"RT";"@SiniOgo:";"Des";"gifles";"se";"perdent";"au";"Senegal";"!";"Un";"seul";"conseil";"prenez";"des";"cours";"de";"self";"défense";"!";"Inscrivez";"vos";"petites";"sœurs";"et";"vos";"fille…"
"Mon Mar 12 14:54:38 CET 2018";"@SunuBuzz Sn";"New";"post:";"Aliou";"Cissé:";"«";"J’ai";"discuté";"avec";"Ferland";"Mendy";"d’une";"possibilité";"de";"jouer";"pour";"le";"Sénégal";"»";"https://t.co/VTxPPkDUJU"
"Mon Mar 12 14:54:15 CET 2018";"@Emmanuel Amunala";"RT";"@oumar_khassoum:";"Hell";"yeah";"🇸🇳🇸🇳🇸🇳";"Senegal";"is";"Bae😜";"#FinePeoplefromSenegal";"";"#FinePeoplefromAfrica";"https://t.co/b3drwboodR"
"Mon Mar 12 14:53:56 CET 2018";"@Boy Next Door 🙎🏾‍♂️";"Senegal";"win";"this";"contest";"❤️❤️";"https://t.co/wvl4sUUl3z"
"Mon Mar 12 14:53:41 CET 2018";"@Maricab";"Sénégal";"-";"Vidéo:";"Professeur";"Songué";"Diouf";"aux";"femmes";"violées";"« Vous";"faites";"tout";"pour";"que";"nous";"vous";"violons »";"https://t.co/FN8QiF4gCX";"via";"@YouTube";"Les";"gens";"autour";"👀";"👀";"👀";"#cultureduviol";"#rapeCulture"
"Mon Mar 12 14:53:31 CET 2018";"@fadel diagne";"RT";"@GalsenHistory:";"Le";""Talatay";"Nder"";"c'etait";"le";"Mardi";"07";"mars";"1820,";"à";"Nder,";"capitale";"du";"Royaume";"du";"Waalo.Ce";"jour";"là,";"la";"Linguère";"Fatim";"Yama…"
"Mon Mar 12 14:53:28 CET 2018";"@Ati Randolph";"RT";"@atrandolph:";"#Togo";"#AshRévolution";"#Direct";"#Live";"#Grève";"Générale";"dans";"toute";"la";"Fonction";"Publique";"!";"Peuple";"Togolais";"tous";"dans";"la";"rue";"et";"su…"
"Mon Mar 12 14:53:17 CET 2018";"@el sarguito";"@pfl1976";"@PensadorZarolho";"Já";"passei";"as";"passas";"do";"Algarve";"ali...";"burrei";"a";"cuequinha";"toda"
"Mon Mar 12 14:53:05 CET 2018";"@Ati Randolph";"RT";"@atrandolph:";"#Togo:";"#URGENT";"deux";"#étudiants";"du";"#frontCitoyen";"#TogoDebout";"arrêtés";"par";"les";"sbires";"du";"#filsDepute";"#Gnassingbé";"";"https://t.co…"
"Mon Mar 12 14:52:47 CET 2018";"@Sassouman";"RT";"@SySeynabou:";"J'invite";"mes";"amis,chercheurs";"ou";"pas,";"qui";"se";"sentent";"concernés";"de";"constituer";"une";"équipe";"pluridisciplinaire";"et";"faire";"1";"étude…"
"Mon Mar 12 14:52:46 CET 2018";"@Donbesh";"RT";"@y___yvss:";"Booba";"interdit";"de";"Lyon";"par";"Bassem,";"interdit";"de";"Senegal";"par";"Alpha,";"interdit";"de";"Comores";"par";"Rohff,";"interdit";"de";"thaïlande";"par";"Se…"
"Mon Mar 12 14:52:28 CET 2018";"@Collateral Beauty";"Éduquez";"vos";"enfants";"correctement.";"Les";"femmes";"parlez(";"é.d.u.q.u.e.z";"les)";"à";"vos";"maris,";"à";"vos";"";"frères";"et";"vos";"cousins.";"On";"en";"a";"marre";"de";"ces";"hommes";"qui";"pensent";"que";"violer";"est";"normal";"ou";"excusable.";"#Senegal"
"Mon Mar 12 14:52:03 CET 2018";"@march24💓";"Dang";"can";"I";"do";"a";"fine";"people";"from";"Senegal";"or";"I";"don’t";"qualify?😂"
"Mon Mar 12 14:51:57 CET 2018";"@Gatabazi JMV";"RT";"@abillen2:";"Le";"Président";"Paul";"#Kagame";"mobilise";"le";"secteur";"privé";"pour";"le";"financement";"de";"l'énergie";"solaire";"(New";"Delhi";"–";"#Inde).";"#Rwanda";"#Ma…"
"Mon Mar 12 14:51:44 CET 2018";"@Diaby Mohamed";"RT";"@SySeynabou:";"J'invite";"mes";"amis,chercheurs";"ou";"pas,";"qui";"se";"sentent";"concernés";"de";"constituer";"une";"équipe";"pluridisciplinaire";"et";"faire";"1";"étude…"
"Mon Mar 12 14:51:29 CET 2018";"@SeneNews";"Urgent-Karang";":";"les";"élèves";"brûlent";"leurs";"blouses";"devant";"l’administration";"#kebetu";"#senegal";"https://t.co/eJRWDjqUgJ";"https://t.co/wUNhVKdPl6"
"Mon Mar 12 14:51:01 CET 2018";"@Todo Sobre Camisetas";"@PabloEstebanCS";"ahí";"ya";"es";"falla";"de";"la";"federación";"de";"Senegal.";"Qué";"falla";"ver";"tantas";"camisetas";"desactualizadas."
"Mon Mar 12 14:50:45 CET 2018";"@DoroFineGirl";"RT";"@SiniOgo:";"Des";"gifles";"se";"perdent";"au";"Senegal";"!";"Un";"seul";"conseil";"prenez";"des";"cours";"de";"self";"défense";"!";"Inscrivez";"vos";"petites";"sœurs";"et";"vos";"fille…"
"Mon Mar 12 14:49:59 CET 2018";"@✝ Contre Яévolution";"RT";"@HRyssen:";"Au";"#Sénégal,";"visiblement,";"une";"bonne";"parti";"du";"commerce";"et";"de";"l'industrie";"sont";"liés";"à";"l'Etat";"hébreu";":";"pétrole,";"engrais,";"pesticid…"
"Mon Mar 12 14:49:35 CET 2018";"@succes | losses";"RT";"@y___yvss:";"Booba";"interdit";"de";"Lyon";"par";"Bassem,";"interdit";"de";"Senegal";"par";"Alpha,";"interdit";"de";"Comores";"par";"Rohff,";"interdit";"de";"thaïlande";"par";"Se…"
"Mon Mar 12 14:49:32 CET 2018";"@TheRealNaala. 🥀";"RT";"@shadyfool:";"Mais";"lui";"là";"il";"est";"caché";"où";"dans";"le";"Sénégal";"?";"https://t.co/yFvl7IiRaq"
"Mon Mar 12 14:49:17 CET 2018";"@Nicolas II";"RT";"@HRyssen:";"Au";"#Sénégal,";"visiblement,";"une";"bonne";"parti";"du";"commerce";"et";"de";"l'industrie";"sont";"liés";"à";"l'Etat";"hébreu";":";"pétrole,";"engrais,";"pesticid…"
"Mon Mar 12 14:49:12 CET 2018";"@Angel⚜️";"N’ayant";"pas";"toute";"ma";"tête";"actuellement,";"une";"bonne";"réflexion";"serait";"un";"peu";"difficile.";"Mais,";"je";"pense";"que";"nous";"avons";"de";"fausses";"opinions,";"des";"réalités";"mensongères";"sur";"le";"mariage";"au";"Sénégal.";"https://t.co/r9HlGZknu0"
"Mon Mar 12 14:48:57 CET 2018";"@Tom Huang";"RT";"@TheDIHC:";"Set";"sail";"to";"Senegal";"with";"Author";"and";"Journalist";"Anna";"Badkhen.";"#flashsale";"";"";"Tuesday,";"March";"13,";"6:30";"pm";"6:00";"pm";"reception";"https:/…"
"Mon Mar 12 14:48:36 CET 2018";"@ibrahim toure";"@SAVE_DAKAR";"Loool...";"C";""la";"senegal";"emergent"";"";"Khadim";"Samb"
"Mon Mar 12 14:48:08 CET 2018";"@seemedeh";"RT";"@LACMA:";"Maïmouna";"Guerresi";"is";"an";"Italian-born";"artist";"who";"converted";"to";"Islam,";"joining";"a";"Sufi";"community";"in";"Senegal";"in";"the";"early";"1990s.";"She…"
"Mon Mar 12 14:47:40 CET 2018";"@IAM A JEADER";"Le";"Super";"Women";"Leadership";"Conference";"2018";"de";"JEADER";"SENEGAL,";"ce";"sera";"ce";"Samedi";"17";"au";"Novotel";"sous";"le";"thème";"de";"la";"Trans'Mission";"!";"Réservez";"votre";"place";"!";"https://t.co/iJriKdI4O5";"@Eventbrite";"@NatyMbaye";"@mamouchkadiop";"@KhadidiatouFSAM";"@mafantadiallo";"@NdyeAbsaGningue";"@PapaCheikhFall2"
"Mon Mar 12 14:47:36 CET 2018";"@Sait Matty Jaw";"RT";"@BarrowPresident:";"We";"belief";"in";"strengthening";"bilateral";"ties";"for";"the";"socio-economic";"and";"political";"benefits";"of";"our";"people.";"";"I";"am";"honoured…"
"Mon Mar 12 14:47:22 CET 2018";"@C.N.I.D.";"Avis";"de";"Recrutement";"d’un(e)";"Chargé(e)";"de";"Programme";"Protection";"de";"l'enfance";"";"Lieu";"d’affectation:";"Bureau";"de";"Pays";"Dakar";"Grade";":";"NOB";"Date";"limite";"de";"soumission:";"23";"Mars";"2018";"Soumettez";"votre";"candidature";"en";"allant";"sur";":";"https://t.co/D75hzjEQr2"
"Mon Mar 12 14:47:19 CET 2018";"@MiLK ®";"RT";"@RicaSenegal:";"Disponible";"Au";"senegal";"https://t.co/YJOB4PBTUp"
"Mon Mar 12 14:47:12 CET 2018";"@WAKANDA";"J’ai";"pas";"regarder";"la";"vidéo";"du";"gars";"là";"dans";"Jakarlo,";"je";"peux";"juste";"pas.";"Oh";"mon";"Senegal...."
